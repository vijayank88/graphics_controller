magic
tech sky130B
magscale 1 2
timestamp 1661955789
<< obsli1 >>
rect 1104 2159 137632 138737
<< obsm1 >>
rect 14 1776 138538 139188
<< metal2 >>
rect 662 140141 718 140941
rect 3882 140141 3938 140941
rect 6458 140141 6514 140941
rect 9678 140141 9734 140941
rect 12254 140141 12310 140941
rect 15474 140141 15530 140941
rect 18694 140141 18750 140941
rect 21270 140141 21326 140941
rect 24490 140141 24546 140941
rect 27066 140141 27122 140941
rect 30286 140141 30342 140941
rect 32862 140141 32918 140941
rect 36082 140141 36138 140941
rect 38658 140141 38714 140941
rect 41878 140141 41934 140941
rect 45098 140141 45154 140941
rect 47674 140141 47730 140941
rect 50894 140141 50950 140941
rect 53470 140141 53526 140941
rect 56690 140141 56746 140941
rect 59266 140141 59322 140941
rect 62486 140141 62542 140941
rect 65706 140141 65762 140941
rect 68282 140141 68338 140941
rect 71502 140141 71558 140941
rect 74078 140141 74134 140941
rect 77298 140141 77354 140941
rect 79874 140141 79930 140941
rect 83094 140141 83150 140941
rect 85670 140141 85726 140941
rect 88890 140141 88946 140941
rect 92110 140141 92166 140941
rect 94686 140141 94742 140941
rect 97906 140141 97962 140941
rect 100482 140141 100538 140941
rect 103702 140141 103758 140941
rect 106278 140141 106334 140941
rect 109498 140141 109554 140941
rect 112074 140141 112130 140941
rect 115294 140141 115350 140941
rect 118514 140141 118570 140941
rect 121090 140141 121146 140941
rect 124310 140141 124366 140941
rect 126886 140141 126942 140941
rect 130106 140141 130162 140941
rect 132682 140141 132738 140941
rect 135902 140141 135958 140941
rect 138478 140141 138534 140941
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 8390 0 8446 800
rect 11610 0 11666 800
rect 14186 0 14242 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 23202 0 23258 800
rect 26422 0 26478 800
rect 28998 0 29054 800
rect 32218 0 32274 800
rect 34794 0 34850 800
rect 38014 0 38070 800
rect 40590 0 40646 800
rect 43810 0 43866 800
rect 46386 0 46442 800
rect 49606 0 49662 800
rect 52826 0 52882 800
rect 55402 0 55458 800
rect 58622 0 58678 800
rect 61198 0 61254 800
rect 64418 0 64474 800
rect 66994 0 67050 800
rect 70214 0 70270 800
rect 72790 0 72846 800
rect 76010 0 76066 800
rect 79230 0 79286 800
rect 81806 0 81862 800
rect 85026 0 85082 800
rect 87602 0 87658 800
rect 90822 0 90878 800
rect 93398 0 93454 800
rect 96618 0 96674 800
rect 99838 0 99894 800
rect 102414 0 102470 800
rect 105634 0 105690 800
rect 108210 0 108266 800
rect 111430 0 111486 800
rect 114006 0 114062 800
rect 117226 0 117282 800
rect 119802 0 119858 800
rect 123022 0 123078 800
rect 126242 0 126298 800
rect 128818 0 128874 800
rect 132038 0 132094 800
rect 134614 0 134670 800
rect 137834 0 137890 800
<< obsm2 >>
rect 20 140085 606 140298
rect 774 140085 3826 140298
rect 3994 140085 6402 140298
rect 6570 140085 9622 140298
rect 9790 140085 12198 140298
rect 12366 140085 15418 140298
rect 15586 140085 18638 140298
rect 18806 140085 21214 140298
rect 21382 140085 24434 140298
rect 24602 140085 27010 140298
rect 27178 140085 30230 140298
rect 30398 140085 32806 140298
rect 32974 140085 36026 140298
rect 36194 140085 38602 140298
rect 38770 140085 41822 140298
rect 41990 140085 45042 140298
rect 45210 140085 47618 140298
rect 47786 140085 50838 140298
rect 51006 140085 53414 140298
rect 53582 140085 56634 140298
rect 56802 140085 59210 140298
rect 59378 140085 62430 140298
rect 62598 140085 65650 140298
rect 65818 140085 68226 140298
rect 68394 140085 71446 140298
rect 71614 140085 74022 140298
rect 74190 140085 77242 140298
rect 77410 140085 79818 140298
rect 79986 140085 83038 140298
rect 83206 140085 85614 140298
rect 85782 140085 88834 140298
rect 89002 140085 92054 140298
rect 92222 140085 94630 140298
rect 94798 140085 97850 140298
rect 98018 140085 100426 140298
rect 100594 140085 103646 140298
rect 103814 140085 106222 140298
rect 106390 140085 109442 140298
rect 109610 140085 112018 140298
rect 112186 140085 115238 140298
rect 115406 140085 118458 140298
rect 118626 140085 121034 140298
rect 121202 140085 124254 140298
rect 124422 140085 126830 140298
rect 126998 140085 130050 140298
rect 130218 140085 132626 140298
rect 132794 140085 135846 140298
rect 136014 140085 138422 140298
rect 20 856 138532 140085
rect 130 800 2538 856
rect 2706 800 5758 856
rect 5926 800 8334 856
rect 8502 800 11554 856
rect 11722 800 14130 856
rect 14298 800 17350 856
rect 17518 800 19926 856
rect 20094 800 23146 856
rect 23314 800 26366 856
rect 26534 800 28942 856
rect 29110 800 32162 856
rect 32330 800 34738 856
rect 34906 800 37958 856
rect 38126 800 40534 856
rect 40702 800 43754 856
rect 43922 800 46330 856
rect 46498 800 49550 856
rect 49718 800 52770 856
rect 52938 800 55346 856
rect 55514 800 58566 856
rect 58734 800 61142 856
rect 61310 800 64362 856
rect 64530 800 66938 856
rect 67106 800 70158 856
rect 70326 800 72734 856
rect 72902 800 75954 856
rect 76122 800 79174 856
rect 79342 800 81750 856
rect 81918 800 84970 856
rect 85138 800 87546 856
rect 87714 800 90766 856
rect 90934 800 93342 856
rect 93510 800 96562 856
rect 96730 800 99782 856
rect 99950 800 102358 856
rect 102526 800 105578 856
rect 105746 800 108154 856
rect 108322 800 111374 856
rect 111542 800 113950 856
rect 114118 800 117170 856
rect 117338 800 119746 856
rect 119914 800 122966 856
rect 123134 800 126186 856
rect 126354 800 128762 856
rect 128930 800 131982 856
rect 132150 800 134558 856
rect 134726 800 137778 856
rect 137946 800 138532 856
<< metal3 >>
rect 0 139408 800 139528
rect 137997 138048 138797 138168
rect 0 136008 800 136128
rect 137997 134648 138797 134768
rect 0 133288 800 133408
rect 137997 131928 138797 132048
rect 0 129888 800 130008
rect 137997 128528 138797 128648
rect 0 126488 800 126608
rect 137997 125808 138797 125928
rect 0 123768 800 123888
rect 137997 122408 138797 122528
rect 0 120368 800 120488
rect 137997 119688 138797 119808
rect 0 117648 800 117768
rect 137997 116288 138797 116408
rect 0 114248 800 114368
rect 137997 112888 138797 113008
rect 0 111528 800 111648
rect 137997 110168 138797 110288
rect 0 108128 800 108248
rect 137997 106768 138797 106888
rect 0 105408 800 105528
rect 137997 104048 138797 104168
rect 0 102008 800 102128
rect 137997 100648 138797 100768
rect 0 98608 800 98728
rect 137997 97928 138797 98048
rect 0 95888 800 96008
rect 137997 94528 138797 94648
rect 0 92488 800 92608
rect 137997 91808 138797 91928
rect 0 89768 800 89888
rect 137997 88408 138797 88528
rect 0 86368 800 86488
rect 137997 85008 138797 85128
rect 0 83648 800 83768
rect 137997 82288 138797 82408
rect 0 80248 800 80368
rect 137997 78888 138797 79008
rect 0 76848 800 76968
rect 137997 76168 138797 76288
rect 0 74128 800 74248
rect 137997 72768 138797 72888
rect 0 70728 800 70848
rect 137997 70048 138797 70168
rect 0 68008 800 68128
rect 137997 66648 138797 66768
rect 0 64608 800 64728
rect 137997 63928 138797 64048
rect 0 61888 800 62008
rect 137997 60528 138797 60648
rect 0 58488 800 58608
rect 137997 57128 138797 57248
rect 0 55768 800 55888
rect 137997 54408 138797 54528
rect 0 52368 800 52488
rect 137997 51008 138797 51128
rect 0 48968 800 49088
rect 137997 48288 138797 48408
rect 0 46248 800 46368
rect 137997 44888 138797 45008
rect 0 42848 800 42968
rect 137997 42168 138797 42288
rect 0 40128 800 40248
rect 137997 38768 138797 38888
rect 0 36728 800 36848
rect 137997 35368 138797 35488
rect 0 34008 800 34128
rect 137997 32648 138797 32768
rect 0 30608 800 30728
rect 137997 29248 138797 29368
rect 0 27888 800 28008
rect 137997 26528 138797 26648
rect 0 24488 800 24608
rect 137997 23128 138797 23248
rect 0 21088 800 21208
rect 137997 20408 138797 20528
rect 0 18368 800 18488
rect 137997 17008 138797 17128
rect 0 14968 800 15088
rect 137997 14288 138797 14408
rect 0 12248 800 12368
rect 137997 10888 138797 11008
rect 0 8848 800 8968
rect 137997 7488 138797 7608
rect 0 6128 800 6248
rect 137997 4768 138797 4888
rect 0 2728 800 2848
rect 137997 1368 138797 1488
<< obsm3 >>
rect 880 139328 137997 139501
rect 800 138248 137997 139328
rect 800 137968 137917 138248
rect 800 136208 137997 137968
rect 880 135928 137997 136208
rect 800 134848 137997 135928
rect 800 134568 137917 134848
rect 800 133488 137997 134568
rect 880 133208 137997 133488
rect 800 132128 137997 133208
rect 800 131848 137917 132128
rect 800 130088 137997 131848
rect 880 129808 137997 130088
rect 800 128728 137997 129808
rect 800 128448 137917 128728
rect 800 126688 137997 128448
rect 880 126408 137997 126688
rect 800 126008 137997 126408
rect 800 125728 137917 126008
rect 800 123968 137997 125728
rect 880 123688 137997 123968
rect 800 122608 137997 123688
rect 800 122328 137917 122608
rect 800 120568 137997 122328
rect 880 120288 137997 120568
rect 800 119888 137997 120288
rect 800 119608 137917 119888
rect 800 117848 137997 119608
rect 880 117568 137997 117848
rect 800 116488 137997 117568
rect 800 116208 137917 116488
rect 800 114448 137997 116208
rect 880 114168 137997 114448
rect 800 113088 137997 114168
rect 800 112808 137917 113088
rect 800 111728 137997 112808
rect 880 111448 137997 111728
rect 800 110368 137997 111448
rect 800 110088 137917 110368
rect 800 108328 137997 110088
rect 880 108048 137997 108328
rect 800 106968 137997 108048
rect 800 106688 137917 106968
rect 800 105608 137997 106688
rect 880 105328 137997 105608
rect 800 104248 137997 105328
rect 800 103968 137917 104248
rect 800 102208 137997 103968
rect 880 101928 137997 102208
rect 800 100848 137997 101928
rect 800 100568 137917 100848
rect 800 98808 137997 100568
rect 880 98528 137997 98808
rect 800 98128 137997 98528
rect 800 97848 137917 98128
rect 800 96088 137997 97848
rect 880 95808 137997 96088
rect 800 94728 137997 95808
rect 800 94448 137917 94728
rect 800 92688 137997 94448
rect 880 92408 137997 92688
rect 800 92008 137997 92408
rect 800 91728 137917 92008
rect 800 89968 137997 91728
rect 880 89688 137997 89968
rect 800 88608 137997 89688
rect 800 88328 137917 88608
rect 800 86568 137997 88328
rect 880 86288 137997 86568
rect 800 85208 137997 86288
rect 800 84928 137917 85208
rect 800 83848 137997 84928
rect 880 83568 137997 83848
rect 800 82488 137997 83568
rect 800 82208 137917 82488
rect 800 80448 137997 82208
rect 880 80168 137997 80448
rect 800 79088 137997 80168
rect 800 78808 137917 79088
rect 800 77048 137997 78808
rect 880 76768 137997 77048
rect 800 76368 137997 76768
rect 800 76088 137917 76368
rect 800 74328 137997 76088
rect 880 74048 137997 74328
rect 800 72968 137997 74048
rect 800 72688 137917 72968
rect 800 70928 137997 72688
rect 880 70648 137997 70928
rect 800 70248 137997 70648
rect 800 69968 137917 70248
rect 800 68208 137997 69968
rect 880 67928 137997 68208
rect 800 66848 137997 67928
rect 800 66568 137917 66848
rect 800 64808 137997 66568
rect 880 64528 137997 64808
rect 800 64128 137997 64528
rect 800 63848 137917 64128
rect 800 62088 137997 63848
rect 880 61808 137997 62088
rect 800 60728 137997 61808
rect 800 60448 137917 60728
rect 800 58688 137997 60448
rect 880 58408 137997 58688
rect 800 57328 137997 58408
rect 800 57048 137917 57328
rect 800 55968 137997 57048
rect 880 55688 137997 55968
rect 800 54608 137997 55688
rect 800 54328 137917 54608
rect 800 52568 137997 54328
rect 880 52288 137997 52568
rect 800 51208 137997 52288
rect 800 50928 137917 51208
rect 800 49168 137997 50928
rect 880 48888 137997 49168
rect 800 48488 137997 48888
rect 800 48208 137917 48488
rect 800 46448 137997 48208
rect 880 46168 137997 46448
rect 800 45088 137997 46168
rect 800 44808 137917 45088
rect 800 43048 137997 44808
rect 880 42768 137997 43048
rect 800 42368 137997 42768
rect 800 42088 137917 42368
rect 800 40328 137997 42088
rect 880 40048 137997 40328
rect 800 38968 137997 40048
rect 800 38688 137917 38968
rect 800 36928 137997 38688
rect 880 36648 137997 36928
rect 800 35568 137997 36648
rect 800 35288 137917 35568
rect 800 34208 137997 35288
rect 880 33928 137997 34208
rect 800 32848 137997 33928
rect 800 32568 137917 32848
rect 800 30808 137997 32568
rect 880 30528 137997 30808
rect 800 29448 137997 30528
rect 800 29168 137917 29448
rect 800 28088 137997 29168
rect 880 27808 137997 28088
rect 800 26728 137997 27808
rect 800 26448 137917 26728
rect 800 24688 137997 26448
rect 880 24408 137997 24688
rect 800 23328 137997 24408
rect 800 23048 137917 23328
rect 800 21288 137997 23048
rect 880 21008 137997 21288
rect 800 20608 137997 21008
rect 800 20328 137917 20608
rect 800 18568 137997 20328
rect 880 18288 137997 18568
rect 800 17208 137997 18288
rect 800 16928 137917 17208
rect 800 15168 137997 16928
rect 880 14888 137997 15168
rect 800 14488 137997 14888
rect 800 14208 137917 14488
rect 800 12448 137997 14208
rect 880 12168 137997 12448
rect 800 11088 137997 12168
rect 800 10808 137917 11088
rect 800 9048 137997 10808
rect 880 8768 137997 9048
rect 800 7688 137997 8768
rect 800 7408 137917 7688
rect 800 6328 137997 7408
rect 880 6048 137997 6328
rect 800 4968 137997 6048
rect 800 4688 137917 4968
rect 800 2928 137997 4688
rect 880 2648 137997 2928
rect 800 1568 137997 2648
rect 800 1395 137917 1568
<< metal4 >>
rect 4208 2128 4528 138768
rect 19568 2128 19888 138768
rect 34928 2128 35248 138768
rect 50288 2128 50608 138768
rect 65648 2128 65968 138768
rect 81008 2128 81328 138768
rect 96368 2128 96688 138768
rect 111728 2128 112048 138768
rect 127088 2128 127408 138768
<< obsm4 >>
rect 4843 2048 19488 138413
rect 19968 2048 34848 138413
rect 35328 2048 50208 138413
rect 50688 2048 65568 138413
rect 66048 2048 80928 138413
rect 81408 2048 96288 138413
rect 96768 2048 111648 138413
rect 112128 2048 127008 138413
rect 127488 2048 136469 138413
rect 4843 1939 136469 2048
<< labels >>
rlabel metal2 s 66994 0 67050 800 6 dbg_freeze_i
port 1 nsew signal input
rlabel metal3 s 137997 138048 138797 138168 6 irq_gfx_o
port 2 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 lt24_cs_n_o
port 3 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 lt24_d_en_o
port 4 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 lt24_d_i[0]
port 5 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 lt24_d_i[10]
port 6 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 lt24_d_i[11]
port 7 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 lt24_d_i[12]
port 8 nsew signal input
rlabel metal3 s 137997 14288 138797 14408 6 lt24_d_i[13]
port 9 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 lt24_d_i[14]
port 10 nsew signal input
rlabel metal3 s 137997 32648 138797 32768 6 lt24_d_i[15]
port 11 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 lt24_d_i[1]
port 12 nsew signal input
rlabel metal2 s 45098 140141 45154 140941 6 lt24_d_i[2]
port 13 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 lt24_d_i[3]
port 14 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 lt24_d_i[4]
port 15 nsew signal input
rlabel metal2 s 77298 140141 77354 140941 6 lt24_d_i[5]
port 16 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 lt24_d_i[6]
port 17 nsew signal input
rlabel metal2 s 38658 140141 38714 140941 6 lt24_d_i[7]
port 18 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 lt24_d_i[8]
port 19 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 lt24_d_i[9]
port 20 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 lt24_d_o[0]
port 21 nsew signal output
rlabel metal2 s 124310 140141 124366 140941 6 lt24_d_o[10]
port 22 nsew signal output
rlabel metal2 s 74078 140141 74134 140941 6 lt24_d_o[11]
port 23 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 lt24_d_o[12]
port 24 nsew signal output
rlabel metal3 s 137997 35368 138797 35488 6 lt24_d_o[13]
port 25 nsew signal output
rlabel metal2 s 27066 140141 27122 140941 6 lt24_d_o[14]
port 26 nsew signal output
rlabel metal3 s 137997 82288 138797 82408 6 lt24_d_o[15]
port 27 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 lt24_d_o[1]
port 28 nsew signal output
rlabel metal2 s 121090 140141 121146 140941 6 lt24_d_o[2]
port 29 nsew signal output
rlabel metal2 s 85670 140141 85726 140941 6 lt24_d_o[3]
port 30 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 lt24_d_o[4]
port 31 nsew signal output
rlabel metal3 s 137997 119688 138797 119808 6 lt24_d_o[5]
port 32 nsew signal output
rlabel metal3 s 137997 104048 138797 104168 6 lt24_d_o[6]
port 33 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 lt24_d_o[7]
port 34 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 lt24_d_o[8]
port 35 nsew signal output
rlabel metal2 s 41878 140141 41934 140941 6 lt24_d_o[9]
port 36 nsew signal output
rlabel metal3 s 137997 106768 138797 106888 6 lt24_on_o
port 37 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 lt24_rd_n_o
port 38 nsew signal output
rlabel metal3 s 137997 17008 138797 17128 6 lt24_reset_n_o
port 39 nsew signal output
rlabel metal3 s 137997 100648 138797 100768 6 lt24_rs_o
port 40 nsew signal output
rlabel metal3 s 137997 42168 138797 42288 6 lt24_wr_n_o
port 41 nsew signal output
rlabel metal2 s 106278 140141 106334 140941 6 lut_ram_addr_o[0]
port 42 nsew signal output
rlabel metal2 s 103702 140141 103758 140941 6 lut_ram_addr_o[1]
port 43 nsew signal output
rlabel metal3 s 137997 125808 138797 125928 6 lut_ram_addr_o[2]
port 44 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 lut_ram_addr_o[3]
port 45 nsew signal output
rlabel metal2 s 30286 140141 30342 140941 6 lut_ram_addr_o[4]
port 46 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 lut_ram_addr_o[5]
port 47 nsew signal output
rlabel metal3 s 137997 134648 138797 134768 6 lut_ram_addr_o[6]
port 48 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 lut_ram_addr_o[7]
port 49 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 lut_ram_addr_o[8]
port 50 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 lut_ram_cen_o
port 51 nsew signal output
rlabel metal3 s 137997 76168 138797 76288 6 lut_ram_din_o[0]
port 52 nsew signal output
rlabel metal3 s 137997 20408 138797 20528 6 lut_ram_din_o[10]
port 53 nsew signal output
rlabel metal2 s 56690 140141 56746 140941 6 lut_ram_din_o[11]
port 54 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 lut_ram_din_o[12]
port 55 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 lut_ram_din_o[13]
port 56 nsew signal output
rlabel metal2 s 662 140141 718 140941 6 lut_ram_din_o[14]
port 57 nsew signal output
rlabel metal3 s 137997 122408 138797 122528 6 lut_ram_din_o[15]
port 58 nsew signal output
rlabel metal3 s 137997 63928 138797 64048 6 lut_ram_din_o[1]
port 59 nsew signal output
rlabel metal2 s 50894 140141 50950 140941 6 lut_ram_din_o[2]
port 60 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 lut_ram_din_o[3]
port 61 nsew signal output
rlabel metal2 s 109498 140141 109554 140941 6 lut_ram_din_o[4]
port 62 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 lut_ram_din_o[5]
port 63 nsew signal output
rlabel metal2 s 130106 140141 130162 140941 6 lut_ram_din_o[6]
port 64 nsew signal output
rlabel metal3 s 137997 1368 138797 1488 6 lut_ram_din_o[7]
port 65 nsew signal output
rlabel metal2 s 126886 140141 126942 140941 6 lut_ram_din_o[8]
port 66 nsew signal output
rlabel metal3 s 137997 26528 138797 26648 6 lut_ram_din_o[9]
port 67 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 lut_ram_dout_i[0]
port 68 nsew signal input
rlabel metal3 s 137997 57128 138797 57248 6 lut_ram_dout_i[10]
port 69 nsew signal input
rlabel metal2 s 115294 140141 115350 140941 6 lut_ram_dout_i[11]
port 70 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 lut_ram_dout_i[12]
port 71 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 lut_ram_dout_i[13]
port 72 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 lut_ram_dout_i[14]
port 73 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 lut_ram_dout_i[15]
port 74 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 lut_ram_dout_i[1]
port 75 nsew signal input
rlabel metal3 s 137997 70048 138797 70168 6 lut_ram_dout_i[2]
port 76 nsew signal input
rlabel metal2 s 53470 140141 53526 140941 6 lut_ram_dout_i[3]
port 77 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 lut_ram_dout_i[4]
port 78 nsew signal input
rlabel metal2 s 15474 140141 15530 140941 6 lut_ram_dout_i[5]
port 79 nsew signal input
rlabel metal3 s 137997 112888 138797 113008 6 lut_ram_dout_i[6]
port 80 nsew signal input
rlabel metal2 s 6458 140141 6514 140941 6 lut_ram_dout_i[7]
port 81 nsew signal input
rlabel metal2 s 32862 140141 32918 140941 6 lut_ram_dout_i[8]
port 82 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 lut_ram_dout_i[9]
port 83 nsew signal input
rlabel metal2 s 71502 140141 71558 140941 6 lut_ram_wen_o
port 84 nsew signal output
rlabel metal2 s 135902 140141 135958 140941 6 mclk
port 85 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 per_addr_i[0]
port 86 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 per_addr_i[10]
port 87 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 per_addr_i[11]
port 88 nsew signal input
rlabel metal2 s 24490 140141 24546 140941 6 per_addr_i[12]
port 89 nsew signal input
rlabel metal3 s 137997 4768 138797 4888 6 per_addr_i[13]
port 90 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 per_addr_i[1]
port 91 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 per_addr_i[2]
port 92 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 per_addr_i[3]
port 93 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 per_addr_i[4]
port 94 nsew signal input
rlabel metal3 s 137997 72768 138797 72888 6 per_addr_i[5]
port 95 nsew signal input
rlabel metal3 s 137997 48288 138797 48408 6 per_addr_i[6]
port 96 nsew signal input
rlabel metal2 s 118514 140141 118570 140941 6 per_addr_i[7]
port 97 nsew signal input
rlabel metal2 s 88890 140141 88946 140941 6 per_addr_i[8]
port 98 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 per_addr_i[9]
port 99 nsew signal input
rlabel metal3 s 137997 131928 138797 132048 6 per_din_i[0]
port 100 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 per_din_i[10]
port 101 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 per_din_i[11]
port 102 nsew signal input
rlabel metal2 s 47674 140141 47730 140941 6 per_din_i[12]
port 103 nsew signal input
rlabel metal2 s 3882 140141 3938 140941 6 per_din_i[13]
port 104 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 per_din_i[14]
port 105 nsew signal input
rlabel metal2 s 12254 140141 12310 140941 6 per_din_i[15]
port 106 nsew signal input
rlabel metal3 s 137997 78888 138797 79008 6 per_din_i[1]
port 107 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 per_din_i[2]
port 108 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 per_din_i[3]
port 109 nsew signal input
rlabel metal3 s 137997 85008 138797 85128 6 per_din_i[4]
port 110 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 per_din_i[5]
port 111 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 per_din_i[6]
port 112 nsew signal input
rlabel metal2 s 59266 140141 59322 140941 6 per_din_i[7]
port 113 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 per_din_i[8]
port 114 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 per_din_i[9]
port 115 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 per_dout_o[0]
port 116 nsew signal output
rlabel metal3 s 137997 54408 138797 54528 6 per_dout_o[10]
port 117 nsew signal output
rlabel metal2 s 62486 140141 62542 140941 6 per_dout_o[11]
port 118 nsew signal output
rlabel metal2 s 83094 140141 83150 140941 6 per_dout_o[12]
port 119 nsew signal output
rlabel metal2 s 79874 140141 79930 140941 6 per_dout_o[13]
port 120 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 per_dout_o[14]
port 121 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 per_dout_o[15]
port 122 nsew signal output
rlabel metal3 s 137997 23128 138797 23248 6 per_dout_o[1]
port 123 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 per_dout_o[2]
port 124 nsew signal output
rlabel metal3 s 137997 116288 138797 116408 6 per_dout_o[3]
port 125 nsew signal output
rlabel metal3 s 137997 88408 138797 88528 6 per_dout_o[4]
port 126 nsew signal output
rlabel metal2 s 92110 140141 92166 140941 6 per_dout_o[5]
port 127 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 per_dout_o[6]
port 128 nsew signal output
rlabel metal3 s 137997 38768 138797 38888 6 per_dout_o[7]
port 129 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 per_dout_o[8]
port 130 nsew signal output
rlabel metal2 s 36082 140141 36138 140941 6 per_dout_o[9]
port 131 nsew signal output
rlabel metal3 s 137997 60528 138797 60648 6 per_en_i
port 132 nsew signal input
rlabel metal3 s 137997 7488 138797 7608 6 per_we_i[0]
port 133 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 per_we_i[1]
port 134 nsew signal input
rlabel metal3 s 137997 110168 138797 110288 6 puc_rst
port 135 nsew signal input
rlabel metal4 s 4208 2128 4528 138768 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 138768 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 138768 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 138768 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 138768 6 vccd1
port 136 nsew power bidirectional
rlabel metal3 s 0 24488 800 24608 6 vid_ram_addr_o[0]
port 137 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 vid_ram_addr_o[10]
port 138 nsew signal output
rlabel metal3 s 137997 44888 138797 45008 6 vid_ram_addr_o[11]
port 139 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 vid_ram_addr_o[12]
port 140 nsew signal output
rlabel metal3 s 137997 10888 138797 11008 6 vid_ram_addr_o[13]
port 141 nsew signal output
rlabel metal2 s 9678 140141 9734 140941 6 vid_ram_addr_o[14]
port 142 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 vid_ram_addr_o[15]
port 143 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 vid_ram_addr_o[16]
port 144 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 vid_ram_addr_o[1]
port 145 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 vid_ram_addr_o[2]
port 146 nsew signal output
rlabel metal3 s 137997 128528 138797 128648 6 vid_ram_addr_o[3]
port 147 nsew signal output
rlabel metal3 s 137997 91808 138797 91928 6 vid_ram_addr_o[4]
port 148 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 vid_ram_addr_o[5]
port 149 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 vid_ram_addr_o[6]
port 150 nsew signal output
rlabel metal3 s 137997 51008 138797 51128 6 vid_ram_addr_o[7]
port 151 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 vid_ram_addr_o[8]
port 152 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 vid_ram_addr_o[9]
port 153 nsew signal output
rlabel metal2 s 138478 140141 138534 140941 6 vid_ram_cen_o
port 154 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 vid_ram_din_o[0]
port 155 nsew signal output
rlabel metal2 s 132682 140141 132738 140941 6 vid_ram_din_o[10]
port 156 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 vid_ram_din_o[11]
port 157 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 vid_ram_din_o[12]
port 158 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 vid_ram_din_o[13]
port 159 nsew signal output
rlabel metal2 s 18 0 74 800 6 vid_ram_din_o[14]
port 160 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 vid_ram_din_o[15]
port 161 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 vid_ram_din_o[1]
port 162 nsew signal output
rlabel metal2 s 18694 140141 18750 140941 6 vid_ram_din_o[2]
port 163 nsew signal output
rlabel metal2 s 68282 140141 68338 140941 6 vid_ram_din_o[3]
port 164 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 vid_ram_din_o[4]
port 165 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 vid_ram_din_o[5]
port 166 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 vid_ram_din_o[6]
port 167 nsew signal output
rlabel metal2 s 94686 140141 94742 140941 6 vid_ram_din_o[7]
port 168 nsew signal output
rlabel metal2 s 65706 140141 65762 140941 6 vid_ram_din_o[8]
port 169 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 vid_ram_din_o[9]
port 170 nsew signal output
rlabel metal2 s 112074 140141 112130 140941 6 vid_ram_dout_i[0]
port 171 nsew signal input
rlabel metal3 s 137997 29248 138797 29368 6 vid_ram_dout_i[10]
port 172 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 vid_ram_dout_i[11]
port 173 nsew signal input
rlabel metal3 s 137997 97928 138797 98048 6 vid_ram_dout_i[12]
port 174 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 vid_ram_dout_i[13]
port 175 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 vid_ram_dout_i[14]
port 176 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 vid_ram_dout_i[15]
port 177 nsew signal input
rlabel metal3 s 137997 94528 138797 94648 6 vid_ram_dout_i[1]
port 178 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 vid_ram_dout_i[2]
port 179 nsew signal input
rlabel metal2 s 100482 140141 100538 140941 6 vid_ram_dout_i[3]
port 180 nsew signal input
rlabel metal2 s 97906 140141 97962 140941 6 vid_ram_dout_i[4]
port 181 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 vid_ram_dout_i[5]
port 182 nsew signal input
rlabel metal2 s 21270 140141 21326 140941 6 vid_ram_dout_i[6]
port 183 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 vid_ram_dout_i[7]
port 184 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 vid_ram_dout_i[8]
port 185 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 vid_ram_dout_i[9]
port 186 nsew signal input
rlabel metal3 s 137997 66648 138797 66768 6 vid_ram_wen_o
port 187 nsew signal output
rlabel metal4 s 19568 2128 19888 138768 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 138768 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 138768 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 138768 6 vssd1
port 188 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 138797 140941
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 51953344
string GDS_FILE /home/vijayan/CARAVEL_FLOW/graphics_controller/openlane/openGFX430/runs/22_08_31_13_48/results/signoff/openGFX430.magic.gds
string GDS_START 1909540
<< end >>

